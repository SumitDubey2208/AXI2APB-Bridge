//
// File: hvl_top.sv
//
// Generated from Mentor VIP Configurator (20191218)
// Generated using Mentor VIP Library ( 2019.4_4 : 10/19/2020:11:53 )
//
module hvl_top;
    import uvm_pkg::*;
    
    `include "test_packages.svh"
    
    initial
    begin
        run_test();
    end

endmodule: hvl_top
