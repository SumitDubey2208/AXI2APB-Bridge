//
// File: test_packages.svh
//
// Generated from Mentor VIP Configurator (20191218)
// Generated using Mentor VIP Library ( 2019.4_4 : 10/19/2020:11:53 )
//

import top_pkg::*;

// Add other packages here as required
