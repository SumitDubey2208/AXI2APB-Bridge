//
// File: top_pkg.sv
//
// Generated from Mentor VIP Configurator (20191218)
// Generated using Mentor VIP Library ( 2019.4_4 : 10/19/2020:11:53 )
//
package top_pkg;
    import uvm_pkg::*;
    
    `include "uvm_macros.svh"
    
    import addr_map_pkg::*;
    
    import top_params_pkg::*;
    import mvc_pkg::*;
    import mgc_axi4_seq_pkg::*;
    import mgc_apb3_v1_0_pkg::*;
    import mgc_axi4_v1_0_pkg::*;
    
    `include "top_env_config.svh"
    `include "top_env.svh"
    `include "top_vseq_base.svh"
    `include "top_test_base.svh"
    `include "top_example_vseq.svh"
endpackage: top_pkg
